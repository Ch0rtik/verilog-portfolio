`default_nettype none
module siren(
	input bit
			clk,
			ENA,
			reset,
			front_door,
			rear_door,
			window,
	input bit [3:0] keypad,
	output bit alarm_siren,
	output bit is_armed,
	output bit is_wait_delay
);
	parameter delay_val = 100;

	bit start_count;
	bit count_done;
	bit [6:0] delay_cntr = 0;
	
	typedef enum bit [1:0] {disarmed, armed, wait_delay, alarm} fsm_states;
	fsm_states curr_state, next_state;

	bit [2:0] sensors;
	assign sensors = {front_door, rear_door, window};
	
	always_ff @(posedge clk)
		if(ENA) begin
			if(reset)
				curr_state <= disarmed;
			else
				curr_state <= next_state;
		end
	
	always_comb 
		unique case(curr_state)
			disarmed: begin 
				if (keypad == 4'b0011)
					next_state <= armed;
				else
					next_state <= curr_state;
			end
			
			armed: begin
				if (sensors != 3'b000)
					next_state <= wait_delay;
				else if (keypad == 4'b1100)
					next_state <= disarmed;
				else 
					next_state <= curr_state;
			end
			
			wait_delay: begin
				if (count_done == 1'b1)
					next_state <= alarm;
				else if (keypad == 4'b1100)
					next_state <= disarmed;
				else 
					next_state <= curr_state;
			end
			
			alarm: begin
				if (keypad == 4'b1100)
					next_state <= disarmed;
				else
					next_state <= curr_state;
			end
		endcase
		
		always_ff @(posedge clk) begin
			if (ENA) begin
				if (reset) begin
					is_armed 		<= 1'b0;
					is_wait_delay 	<= 1'b0;
					alarm_siren		<= 1'b0;
				end else begin
					is_armed			<= (next_state == armed);
					is_wait_delay	<= (next_state == wait_delay);
					alarm_siren		<= (next_state == alarm);
				end
			end
		end
		assign start_count = ((curr_state == armed) && (sensors != 3'b000));
	
		always @(posedge clk)
			if(ENA) begin
				if (reset) 
					delay_cntr <= 7'b0;
				else if (start_count)
					delay_cntr <= delay_val - 7'b1;
				else if (curr_state != wait_delay)
					delay_cntr <= 7'b0;
				else if (delay_cntr != 0)
					delay_cntr <= delay_cntr - 7'b1;
			end
		
		assign count_done = (delay_cntr == 0);

endmodule
